module udp_wrapper (
    input i_clk,
    input i_clk90,
    input i_rst,
    // input i_rst_n,
    output        udp_rx_valid,
    input         udp_rx_ready,
    output        udp_rx_last,
    output [7:0]  udp_rx_data,
    
    input         udp_tx_hdr_valid,
    output  logic udp_tx_hdr_ready,
    output  logic udp_tx_ready,
    input [7:0]   udp_tx_data,
    input         udp_tx_valid,
    input         udp_tx_last,
    // input  [15:0] udp_tx_length,
    
    output [17:0] led_r,
    output [6:0]  hex0,
    output [6:0]  hex1,
    output [6:0]  hex2,
    output [6:0]  hex3,
    output [6:0]  hex4,
    output [6:0]  hex5,
    output [6:0]  hex6,
    output [6:0]  hex7,

    /*
     * Ethernet: 1000BASE-T RGMII
     */
    input        phy0_rx_clk,
    input  [3:0] phy0_rxd,
    input        phy0_rx_ctl,
    output       phy0_tx_clk,
    output [3:0] phy0_txd,
    output       phy0_tx_ctl,
    output       phy0_reset_n,
    input        phy0_int_n

);

// Ethernet Configuration
parameter [47:0] local_mac   = 48'h02_00_00_00_00_00;
parameter [31:0] local_ip    = {8'd192, 8'd168, 8'd50,  8'd168};
parameter [31:0] dest_ip     = {8'd192, 8'd168, 8'd50,  8'd82};
parameter [31:0] gateway_ip  = {8'd192, 8'd168, 8'd50,  8'd1};
parameter [31:0] subnet_mask = {8'd255, 8'd255, 8'd255, 8'd0};
parameter [15:0] udp_port    = 16'd1234;
parameter [15:0] dest_port   = 16'd8080;

// rst
// logic rst;
// assign rst = ~i_rst_n;
assign phy0_reset_n = ~i_rst;

// AXI between MAC and Ethernet modules
logic [7:0] rx_axis_tdata;
logic rx_axis_tvalid;
logic rx_axis_tready;
logic rx_axis_tlast;
logic rx_axis_tuser;

logic [7:0] tx_axis_tdata;
logic tx_axis_tvalid;
logic tx_axis_tready;
logic tx_axis_tlast;
logic tx_axis_tuser;

// Ethernet frame between Ethernet modules and UDP stack
logic rx_eth_hdr_ready;
logic rx_eth_hdr_valid;
logic [47:0] rx_eth_dest_mac;
logic [47:0] rx_eth_src_mac;
logic [15:0] rx_eth_type;
logic [7:0] rx_eth_payload_axis_tdata;
logic rx_eth_payload_axis_tvalid;
logic rx_eth_payload_axis_tready;
logic rx_eth_payload_axis_tlast;
logic rx_eth_payload_axis_tuser;

logic tx_eth_hdr_ready;
logic tx_eth_hdr_valid;
logic [47:0] tx_eth_dest_mac;
logic [47:0] tx_eth_src_mac;
logic [15:0] tx_eth_type;
logic [7:0] tx_eth_payload_axis_tdata;
logic tx_eth_payload_axis_tvalid;
logic tx_eth_payload_axis_tready;
logic tx_eth_payload_axis_tlast;
logic tx_eth_payload_axis_tuser;

// IP frame connections
logic rx_ip_hdr_valid;
logic rx_ip_hdr_ready;
logic [47:0] rx_ip_eth_dest_mac;
logic [47:0] rx_ip_eth_src_mac;
logic [15:0] rx_ip_eth_type;
logic [3:0] rx_ip_version;
logic [3:0] rx_ip_ihl;
logic [5:0] rx_ip_dscp;
logic [1:0] rx_ip_ecn;
logic [15:0] rx_ip_length;
logic [15:0] rx_ip_identification;
logic [2:0] rx_ip_flags;
logic [12:0] rx_ip_fragment_offset;
logic [7:0] rx_ip_ttl;
logic [7:0] rx_ip_protocol;
logic [15:0] rx_ip_header_checksum;
logic [31:0] rx_ip_source_ip;
logic [31:0] rx_ip_dest_ip;
logic [7:0] rx_ip_payload_axis_tdata;
logic rx_ip_payload_axis_tvalid;
logic rx_ip_payload_axis_tready;
logic rx_ip_payload_axis_tlast;
logic rx_ip_payload_axis_tuser;

logic tx_ip_hdr_valid;
logic tx_ip_hdr_ready;
logic [5:0] tx_ip_dscp;
logic [1:0] tx_ip_ecn;
logic [15:0] tx_ip_length;
logic [7:0] tx_ip_ttl;
logic [7:0] tx_ip_protocol;
logic [31:0] tx_ip_source_ip;
logic [31:0] tx_ip_dest_ip;
logic [7:0] tx_ip_payload_axis_tdata;
logic tx_ip_payload_axis_tvalid;
logic tx_ip_payload_axis_tready;
logic tx_ip_payload_axis_tlast;
logic tx_ip_payload_axis_tuser;

// UDP frame connections
logic rx_udp_hdr_valid;
logic rx_udp_hdr_ready;
logic [47:0] rx_udp_eth_dest_mac;
logic [47:0] rx_udp_eth_src_mac;
logic [15:0] rx_udp_eth_type;
logic [3:0] rx_udp_ip_version;
logic [3:0] rx_udp_ip_ihl;
logic [5:0] rx_udp_ip_dscp;
logic [1:0] rx_udp_ip_ecn;
logic [15:0] rx_udp_ip_length;
logic [15:0] rx_udp_ip_identification;
logic [2:0] rx_udp_ip_flags;
logic [12:0] rx_udp_ip_fragment_offset;
logic [7:0] rx_udp_ip_ttl;
logic [7:0] rx_udp_ip_protocol;
logic [15:0] rx_udp_ip_header_checksum;
logic [31:0] rx_udp_ip_source_ip;
logic [31:0] rx_udp_ip_dest_ip;
logic [15:0] rx_udp_source_port;
logic [15:0] rx_udp_dest_port;
logic [15:0] rx_udp_length;
logic [15:0] rx_udp_checksum;
logic [7:0] rx_udp_payload_axis_tdata;
logic rx_udp_payload_axis_tvalid;
logic rx_udp_payload_axis_tready;
logic rx_udp_payload_axis_tlast;
logic rx_udp_payload_axis_tuser;

logic tx_udp_hdr_valid;
logic tx_udp_hdr_ready;
logic [5:0] tx_udp_ip_dscp;
logic [1:0] tx_udp_ip_ecn;
logic [7:0] tx_udp_ip_ttl;
logic [31:0] tx_udp_ip_source_ip;
logic [31:0] tx_udp_ip_dest_ip;
logic [15:0] tx_udp_source_port;
logic [15:0] tx_udp_dest_port;
logic [15:0] tx_udp_length;
logic [15:0] tx_udp_checksum;
logic [7:0] tx_udp_payload_axis_tdata;
logic tx_udp_payload_axis_tvalid;
logic tx_udp_payload_axis_tready;
logic tx_udp_payload_axis_tlast;
logic tx_udp_payload_axis_tuser;

logic [7:0] rx_fifo_udp_payload_axis_tdata;
logic rx_fifo_udp_payload_axis_tvalid;
logic rx_fifo_udp_payload_axis_tready;
logic rx_fifo_udp_payload_axis_tlast;
logic rx_fifo_udp_payload_axis_tuser;

logic [7:0] tx_fifo_udp_payload_axis_tdata;
logic tx_fifo_udp_payload_axis_tvalid;
logic tx_fifo_udp_payload_axis_tready;
logic tx_fifo_udp_payload_axis_tlast;
logic tx_fifo_udp_payload_axis_tuser;

// IP ports not used
assign rx_ip_hdr_ready = 1;
assign rx_ip_payload_axis_tready = 1;

assign tx_ip_hdr_valid = 0;
assign tx_ip_dscp = 0;
assign tx_ip_ecn = 0;
assign tx_ip_length = 0;
assign tx_ip_ttl = 0;
assign tx_ip_protocol = 0;
assign tx_ip_source_ip = 0;
assign tx_ip_dest_ip = 0;
assign tx_ip_payload_axis_tdata = 0;
assign tx_ip_payload_axis_tvalid = 0;
assign tx_ip_payload_axis_tlast = 0;
assign tx_ip_payload_axis_tuser = 0;

// assign udp_tx_ready
// assign udp_tx_length
// assign udp_rx_valid = tx_fifo_udp_payload_axis_tvalid;
// assign udp_rx_ready = 
// assign udp_rx_last = tx_fifo_udp_payload_axis_tlast;
// assign udp_data_rx = tx_fifo_udp_payload_axis_tdata;
// assign udp_tx_data

logic match_cond;
assign match_cond = rx_udp_dest_port == 1234;
logic no_match;
assign no_match = !match_cond;
logic match_cond_reg = 0;
logic no_match_reg = 0;

always_ff @(posedge i_clk) begin

    if (i_rst) begin
        match_cond_reg <= 0;
        no_match_reg <= 0;
    end else begin
        if (rx_udp_payload_axis_tvalid) begin
            if ((!match_cond_reg && !no_match_reg) ||
                (rx_udp_payload_axis_tvalid && rx_udp_payload_axis_tready && rx_udp_payload_axis_tlast)) begin
                match_cond_reg <= match_cond;
                no_match_reg <= no_match;
            end
        end else begin
            match_cond_reg <= 0;
            no_match_reg <= 0;
        end
    end
end



assign rx_udp_hdr_ready = (tx_eth_hdr_ready && match_cond) || no_match;

// tx data
assign tx_udp_hdr_valid = udp_tx_hdr_valid;
assign udp_tx_hdr_ready = tx_udp_hdr_ready;


assign tx_udp_ip_dscp = 0;
assign tx_udp_ip_ecn = 0;
assign tx_udp_ip_ttl = 64;
assign tx_udp_ip_source_ip = local_ip;
assign tx_udp_ip_dest_ip = dest_ip;
assign tx_udp_source_port = udp_port;
assign tx_udp_dest_port = dest_port;
assign tx_udp_length = 16'd10;
assign tx_udp_checksum = 0;

// output wire
// assign tx_fifo_udp_payload_axis_tready = tx_udp_payload_axis_tready;
// assign tx_udp_payload_axis_tdata = tx_fifo_udp_payload_axis_tdata;
// assign tx_udp_payload_axis_tvalid = tx_fifo_udp_payload_axis_tvalid;
// assign tx_udp_payload_axis_tlast = tx_fifo_udp_payload_axis_tlast;
assign tx_udp_payload_axis_tuser = tx_fifo_udp_payload_axis_tuser;
// loop back
// assign tx_udp_payload_axis_tdata = udp_rx_data;
// assign tx_udp_payload_axis_tvalid = udp_rx_valid && udp_rx_ready;
assign tx_udp_payload_axis_tvalid = udp_tx_valid;
assign tx_udp_payload_axis_tlast = udp_tx_last;
assign tx_udp_payload_axis_tdata = udp_tx_data;
// assign tx_udp_payload_axis_tvalid = udp_tx_valid;
// assign tx_udp_payload_axis_tlast = udp_tx_last;
// assign udp_tx_ready = udp_rx_valid && udp_rx_ready;
assign udp_tx_ready = tx_udp_payload_axis_tready;


assign rx_fifo_udp_payload_axis_tdata = rx_udp_payload_axis_tdata;
assign rx_fifo_udp_payload_axis_tvalid = rx_udp_payload_axis_tvalid && match_cond_reg;
assign rx_udp_payload_axis_tready = (rx_fifo_udp_payload_axis_tready && match_cond_reg) || no_match_reg;
assign rx_fifo_udp_payload_axis_tlast = rx_udp_payload_axis_tlast;
assign rx_fifo_udp_payload_axis_tuser = rx_udp_payload_axis_tuser;

// Place first payload byte onto LEDs
logic valid_last = 0;
logic [17:0] led_reg_r;

assign led_r = led_reg_r;

always_ff @(posedge i_clk) begin
    
    if (udp_rx_valid) begin
        if (!valid_last) begin
            led_reg_r <= udp_rx_data;
            valid_last <= 1'b1;
        end
        if (udp_rx_last) begin
            valid_last <= 1'b0;
        end
    end

    if (i_rst) begin
        led_reg_r <= 0;
    end
end

// place dest IP onto 7 segment displays
logic [31:0] dest_ip_reg = 0;

always @(posedge i_clk) begin
    if (tx_udp_hdr_valid) begin
        dest_ip_reg <= tx_udp_ip_dest_ip;
    end

    if (i_rst) begin
        dest_ip_reg <= 0;
    end
end

hex_display #(
    .INVERT(1)
)
hex_display_0 (
    .in(dest_ip_reg[3:0]),
    .enable(1),
    .out(hex0)
);

hex_display #(
    .INVERT(1)
)
hex_display_1 (
    .in(dest_ip_reg[7:4]),
    .enable(1),
    .out(hex1)
);

hex_display #(
    .INVERT(1)
)
hex_display_2 (
    .in(dest_ip_reg[11:8]),
    .enable(1),
    .out(hex2)
);

hex_display #(
    .INVERT(1)
)
hex_display_3 (
    .in(dest_ip_reg[15:12]),
    .enable(1),
    .out(hex3)
);

hex_display #(
    .INVERT(1)
)
hex_display_4 (
    .in(dest_ip_reg[19:16]),
    .enable(1),
    .out(hex4)
);

hex_display #(
    .INVERT(1)
)
hex_display_5 (
    .in(dest_ip_reg[23:20]),
    .enable(1),
    .out(hex5)
);

hex_display #(
    .INVERT(1)
)
hex_display_6 (
    .in(dest_ip_reg[27:24]),
    .enable(1),
    .out(hex6)
);

hex_display #(
    .INVERT(1)
)
hex_display_7 (
    .in(dest_ip_reg[31:28]),
    .enable(1),
    .out(hex7)
);


eth_mac_1g_rgmii_fifo #(
    .TARGET("ALTERA"),
    .USE_CLK90("TRUE"),
    .ENABLE_PADDING(1),
    .MIN_FRAME_LENGTH(64),
    .TX_FIFO_DEPTH(4096),
    .TX_FRAME_FIFO(1),
    .RX_FIFO_DEPTH(4096),
    .RX_FRAME_FIFO(1)
)
eth_mac_inst (
    .gtx_clk(i_clk),
    .gtx_clk90(i_clk90),
    .gtx_rst(i_rst),
    .logic_clk(i_clk),
    .logic_rst(i_rst),

    .tx_axis_tdata(tx_axis_tdata),
    .tx_axis_tvalid(tx_axis_tvalid),
    .tx_axis_tready(tx_axis_tready),
    .tx_axis_tlast(tx_axis_tlast),
    .tx_axis_tuser(tx_axis_tuser),
    .rx_axis_tdata(rx_axis_tdata),
    .rx_axis_tvalid(rx_axis_tvalid),
    .rx_axis_tready(rx_axis_tready),
    .rx_axis_tlast(rx_axis_tlast),
    .rx_axis_tuser(rx_axis_tuser),

    .rgmii_rx_clk(phy0_rx_clk),
    .rgmii_rxd(phy0_rxd),
    .rgmii_rx_ctl(phy0_rx_ctl),
    .rgmii_tx_clk(phy0_tx_clk),
    .rgmii_txd(phy0_txd),
    .rgmii_tx_ctl(phy0_tx_ctl),
    
    .tx_fifo_overflow(),
    .tx_fifo_bad_frame(),
    .tx_fifo_good_frame(),
    .rx_error_bad_frame(),
    .rx_error_bad_fcs(),
    .rx_fifo_overflow(),
    .rx_fifo_bad_frame(),
    .rx_fifo_good_frame(),
    .speed(),

    .ifg_delay(12)
);

eth_axis_rx eth_axis_rx_inst (
    .clk(i_clk),
    .rst(i_rst),
    // AXI input
    .s_axis_tdata(rx_axis_tdata),
    .s_axis_tvalid(rx_axis_tvalid),
    .s_axis_tready(rx_axis_tready),
    .s_axis_tlast(rx_axis_tlast),
    .s_axis_tuser(rx_axis_tuser),
    // Ethernet frame output
    .m_eth_hdr_valid(rx_eth_hdr_valid),
    .m_eth_hdr_ready(rx_eth_hdr_ready),
    .m_eth_dest_mac(rx_eth_dest_mac),
    .m_eth_src_mac(rx_eth_src_mac),
    .m_eth_type(rx_eth_type),
    .m_eth_payload_axis_tdata(rx_eth_payload_axis_tdata),
    .m_eth_payload_axis_tvalid(rx_eth_payload_axis_tvalid),
    .m_eth_payload_axis_tready(rx_eth_payload_axis_tready),
    .m_eth_payload_axis_tlast(rx_eth_payload_axis_tlast),
    .m_eth_payload_axis_tuser(rx_eth_payload_axis_tuser),
    // Status signals
    .busy(),
    .error_header_early_termination()
);

eth_axis_tx
eth_axis_tx_inst (
    .clk(i_clk),
    .rst(i_rst),
    // Ethernet frame input
    .s_eth_hdr_valid(tx_eth_hdr_valid),
    .s_eth_hdr_ready(tx_eth_hdr_ready),
    .s_eth_dest_mac(tx_eth_dest_mac),
    .s_eth_src_mac(tx_eth_src_mac),
    .s_eth_type(tx_eth_type),
    .s_eth_payload_axis_tdata(tx_eth_payload_axis_tdata),
    .s_eth_payload_axis_tvalid(tx_eth_payload_axis_tvalid),
    .s_eth_payload_axis_tready(tx_eth_payload_axis_tready),
    .s_eth_payload_axis_tlast(tx_eth_payload_axis_tlast),
    .s_eth_payload_axis_tuser(tx_eth_payload_axis_tuser),
    // AXI output
    .m_axis_tdata(tx_axis_tdata),
    .m_axis_tvalid(tx_axis_tvalid),
    .m_axis_tready(tx_axis_tready),
    .m_axis_tlast(tx_axis_tlast),
    .m_axis_tuser(tx_axis_tuser),
    // Status signals
    .busy()
);

udp_complete
udp_complete_inst (
    .clk(i_clk),
    .rst(i_rst),
    // Ethernet frame input
    .s_eth_hdr_valid(rx_eth_hdr_valid),
    .s_eth_hdr_ready(rx_eth_hdr_ready),
    .s_eth_dest_mac(rx_eth_dest_mac),
    .s_eth_src_mac(rx_eth_src_mac),
    .s_eth_type(rx_eth_type),
    .s_eth_payload_axis_tdata(rx_eth_payload_axis_tdata),
    .s_eth_payload_axis_tvalid(rx_eth_payload_axis_tvalid),
    .s_eth_payload_axis_tready(rx_eth_payload_axis_tready),
    .s_eth_payload_axis_tlast(rx_eth_payload_axis_tlast),
    .s_eth_payload_axis_tuser(rx_eth_payload_axis_tuser),
    // Ethernet frame output
    .m_eth_hdr_valid(tx_eth_hdr_valid),
    .m_eth_hdr_ready(tx_eth_hdr_ready),
    .m_eth_dest_mac(tx_eth_dest_mac),
    .m_eth_src_mac(tx_eth_src_mac),
    .m_eth_type(tx_eth_type),
    .m_eth_payload_axis_tdata(tx_eth_payload_axis_tdata),
    .m_eth_payload_axis_tvalid(tx_eth_payload_axis_tvalid),
    .m_eth_payload_axis_tready(tx_eth_payload_axis_tready),
    .m_eth_payload_axis_tlast(tx_eth_payload_axis_tlast),
    .m_eth_payload_axis_tuser(tx_eth_payload_axis_tuser),
    // IP frame input
    .s_ip_hdr_valid(tx_ip_hdr_valid),
    .s_ip_hdr_ready(tx_ip_hdr_ready),
    .s_ip_dscp(tx_ip_dscp),
    .s_ip_ecn(tx_ip_ecn),
    .s_ip_length(tx_ip_length),
    .s_ip_ttl(tx_ip_ttl),
    .s_ip_protocol(tx_ip_protocol),
    .s_ip_source_ip(tx_ip_source_ip),
    .s_ip_dest_ip(tx_ip_dest_ip),
    .s_ip_payload_axis_tdata(tx_ip_payload_axis_tdata),
    .s_ip_payload_axis_tvalid(tx_ip_payload_axis_tvalid),
    .s_ip_payload_axis_tready(tx_ip_payload_axis_tready),
    .s_ip_payload_axis_tlast(tx_ip_payload_axis_tlast),
    .s_ip_payload_axis_tuser(tx_ip_payload_axis_tuser),
    // IP frame output
    .m_ip_hdr_valid(rx_ip_hdr_valid),
    .m_ip_hdr_ready(rx_ip_hdr_ready),
    .m_ip_eth_dest_mac(rx_ip_eth_dest_mac),
    .m_ip_eth_src_mac(rx_ip_eth_src_mac),
    .m_ip_eth_type(rx_ip_eth_type),
    .m_ip_version(rx_ip_version),
    .m_ip_ihl(rx_ip_ihl),
    .m_ip_dscp(rx_ip_dscp),
    .m_ip_ecn(rx_ip_ecn),
    .m_ip_length(rx_ip_length),
    .m_ip_identification(rx_ip_identification),
    .m_ip_flags(rx_ip_flags),
    .m_ip_fragment_offset(rx_ip_fragment_offset),
    .m_ip_ttl(rx_ip_ttl),
    .m_ip_protocol(rx_ip_protocol),
    .m_ip_header_checksum(rx_ip_header_checksum),
    .m_ip_source_ip(rx_ip_source_ip),
    .m_ip_dest_ip(rx_ip_dest_ip),
    .m_ip_payload_axis_tdata(rx_ip_payload_axis_tdata),
    .m_ip_payload_axis_tvalid(rx_ip_payload_axis_tvalid),
    .m_ip_payload_axis_tready(rx_ip_payload_axis_tready),
    .m_ip_payload_axis_tlast(rx_ip_payload_axis_tlast),
    .m_ip_payload_axis_tuser(rx_ip_payload_axis_tuser),
    // UDP frame input
    .s_udp_hdr_valid(tx_udp_hdr_valid),
    .s_udp_hdr_ready(tx_udp_hdr_ready),
    .s_udp_ip_dscp(tx_udp_ip_dscp),
    .s_udp_ip_ecn(tx_udp_ip_ecn),
    .s_udp_ip_ttl(tx_udp_ip_ttl),
    .s_udp_ip_source_ip(tx_udp_ip_source_ip),
    .s_udp_ip_dest_ip(tx_udp_ip_dest_ip),
    .s_udp_source_port(tx_udp_source_port),
    .s_udp_dest_port(tx_udp_dest_port),
    .s_udp_length(tx_udp_length),
    .s_udp_checksum(tx_udp_checksum),
    // loop back here
    .s_udp_payload_axis_tdata(tx_udp_payload_axis_tdata),
    .s_udp_payload_axis_tvalid(tx_udp_payload_axis_tvalid),
    .s_udp_payload_axis_tready(tx_udp_payload_axis_tready),
    .s_udp_payload_axis_tlast(tx_udp_payload_axis_tlast),
    .s_udp_payload_axis_tuser(tx_udp_payload_axis_tuser),
    // UDP frame output
    .m_udp_hdr_valid(rx_udp_hdr_valid),
    .m_udp_hdr_ready(rx_udp_hdr_ready),
    .m_udp_eth_dest_mac(rx_udp_eth_dest_mac),
    .m_udp_eth_src_mac(rx_udp_eth_src_mac),
    .m_udp_eth_type(rx_udp_eth_type),
    .m_udp_ip_version(rx_udp_ip_version),
    .m_udp_ip_ihl(rx_udp_ip_ihl),
    .m_udp_ip_dscp(rx_udp_ip_dscp),
    .m_udp_ip_ecn(rx_udp_ip_ecn),
    .m_udp_ip_length(rx_udp_ip_length),
    .m_udp_ip_identification(rx_udp_ip_identification),
    .m_udp_ip_flags(rx_udp_ip_flags),
    .m_udp_ip_fragment_offset(rx_udp_ip_fragment_offset),
    .m_udp_ip_ttl(rx_udp_ip_ttl),
    .m_udp_ip_protocol(rx_udp_ip_protocol),
    .m_udp_ip_header_checksum(rx_udp_ip_header_checksum),
    .m_udp_ip_source_ip(rx_udp_ip_source_ip),
    .m_udp_ip_dest_ip(rx_udp_ip_dest_ip),
    .m_udp_source_port(rx_udp_source_port),
    .m_udp_dest_port(rx_udp_dest_port),
    .m_udp_length(rx_udp_length),
    .m_udp_checksum(rx_udp_checksum),
    .m_udp_payload_axis_tdata(rx_udp_payload_axis_tdata),
    .m_udp_payload_axis_tvalid(rx_udp_payload_axis_tvalid),
    .m_udp_payload_axis_tready(rx_udp_payload_axis_tready),
    .m_udp_payload_axis_tlast(rx_udp_payload_axis_tlast),
    .m_udp_payload_axis_tuser(rx_udp_payload_axis_tuser),
    // Status signals
    .ip_rx_busy(),
    .ip_tx_busy(),
    .udp_rx_busy(),
    .udp_tx_busy(),
    .ip_rx_error_header_early_termination(),
    .ip_rx_error_payload_early_termination(),
    .ip_rx_error_invalid_header(),
    .ip_rx_error_invalid_checksum(),
    .ip_tx_error_payload_early_termination(),
    .ip_tx_error_arp_failed(),
    .udp_rx_error_header_early_termination(),
    .udp_rx_error_payload_early_termination(),
    .udp_tx_error_payload_early_termination(),
    // Configuration
    .local_mac(local_mac),
    .local_ip(local_ip),
    .gateway_ip(gateway_ip),
    .subnet_mask(subnet_mask),
    .clear_arp_cache(0)
);

axis_fifo #(
    .DEPTH(8192),
    .DATA_WIDTH(8),
    .KEEP_ENABLE(0),
    .ID_ENABLE(0),
    .DEST_ENABLE(0),
    .USER_ENABLE(1),
    .USER_WIDTH(1),
    .FRAME_FIFO(0)
)
udp_payload_fifo (
    .clk(i_clk),
    .rst(i_rst),

    // AXI input
    .s_axis_tdata(rx_fifo_udp_payload_axis_tdata),
    .s_axis_tkeep(0),
    .s_axis_tvalid(rx_fifo_udp_payload_axis_tvalid),
    .s_axis_tready(rx_fifo_udp_payload_axis_tready),
    .s_axis_tlast(rx_fifo_udp_payload_axis_tlast),
    .s_axis_tid(0),
    .s_axis_tdest(0),
    .s_axis_tuser(rx_fifo_udp_payload_axis_tuser),

    // AXI output
    .m_axis_tdata(udp_rx_data),
    .m_axis_tkeep(),
    .m_axis_tvalid(udp_rx_valid),
    .m_axis_tready(udp_rx_ready),
    .m_axis_tlast(udp_rx_last),
    .m_axis_tid(),
    .m_axis_tdest(),
    .m_axis_tuser(tx_fifo_udp_payload_axis_tuser),

    // Status
    .status_overflow(),
    .status_bad_frame(),
    .status_good_frame()
);


endmodule