module receiver (
    input 
);
    
endmodule